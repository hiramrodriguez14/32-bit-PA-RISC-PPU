module mux32x5 (
    input [31:0] R0, R1, R2, R3, R4, R5, R6, R7, R8, R9,
                 R10, R11, R12, R13, R14, R15, R16, R17, R18, R19,
                 R20, R21, R22, R23, R24, R25, R26, R27, R28, R29,
                 R30, R31,  
    input [4:0] S,          // 5-bit selector
    output wire [31:0] N    // Selected output
);

    assign N = (S == 5'd0)  ? R0  :
               (S == 5'd1)  ? R1  :
               (S == 5'd2)  ? R2  :
               (S == 5'd3)  ? R3  :
               (S == 5'd4)  ? R4  :
               (S == 5'd5)  ? R5  :
               (S == 5'd6)  ? R6  :
               (S == 5'd7)  ? R7  :
               (S == 5'd8)  ? R8  :
               (S == 5'd9)  ? R9  :
               (S == 5'd10) ? R10 :
               (S == 5'd11) ? R11 :
               (S == 5'd12) ? R12 :
               (S == 5'd13) ? R13 :
               (S == 5'd14) ? R14 :
               (S == 5'd15) ? R15 :
               (S == 5'd16) ? R16 :
               (S == 5'd17) ? R17 :
               (S == 5'd18) ? R18 :
               (S == 5'd19) ? R19 :
               (S == 5'd20) ? R20 :
               (S == 5'd21) ? R21 :
               (S == 5'd22) ? R22 :
               (S == 5'd23) ? R23 :
               (S == 5'd24) ? R24 :
               (S == 5'd25) ? R25 :
               (S == 5'd26) ? R26 :
               (S == 5'd27) ? R27 :
               (S == 5'd28) ? R28 :
               (S == 5'd29) ? R29 :
               (S == 5'd30) ? R30 :
               (S == 5'd31) ? R31 :
                             32'b0;
endmodule
